module data_memory #(
    parameter ADDRESS_WIDTH = 32,
              DATA_WIDTH = 32
)(
    //diagram specifies wr_en_i only so will always be reading/ writing. No re_en_i.
    //also specifies one address in
    input logic clk_i,
    input logic wr_en_i,
    input logic [ADDRESS_WIDTH-1:0] addr_i,
    input logic [DATA_WIDTH-1:0] data_i,
    output logic [DATA_WIDTH-1:0] data_o
);

logic [7:0] ram_array [131071-1:0];

initial begin
    for (int i = 0; i < 131072; i++) begin
        ram_array[i]=8'b0;
    end
    $readmemh("sine.mem", ram_array, "h10000");
end

always_ff @(posedge clk_i) begin
    if (wr_en_i == 1'b1)
        ram_array[addr_i] <= data_i;
    else
        // output is synchronous
        data_o <= ram_array[addr_i];
end

endmodule
